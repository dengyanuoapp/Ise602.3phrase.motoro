module m3_powerAndSpeedCalc (
    
    clkI,
    nRstI
)
input   wire                m3startI;	
input   wire                m3forceStopI;	 
input   wire                m3invRotateI;	 
input   wire                m3freqINCi	;
input   wire                m3freqDECi	;
input   wire                m3powerINCi	;
input   wire                m3powerDECi	;

input wire                  clkI       ;
input wire                  nRstI      ;
